Library IEEE;
Use IEEE.STD_LOGIC_1164.ALL;
Use IEEE.STD_LOGIC_ARITH.ALL;
Use IEEE.STD_LOGIC_UNSIGNED.ALL;

Entity half_add is
	Port(A : in std_logic;
		  B : in std_logic;
		  C : out std_logic;
		  S : out std_logic);
End half_add;

Architecture Behavioral of half_add is
Begin
	C <= A and B;
	S <= A xor B;
End Behavioral;